module ALU(read_data_1,read_data_2,ALUcontrol,ALUresult);
  
  input read_data_1[4:0],read_data_2[4:0],ALUcontrol[4:0];
  output ALUresult